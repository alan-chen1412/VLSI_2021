//================================================
// Auther:      Chang Wan-Yun (Claire)            
// Filename:    AXI.sv                            
// Description: Top module of AXI                  
// Version:     1.0 
//================================================
`include "AXI_master_p.sv"
`include "AXI_slave_p.sv"
`include "Arbiter.sv"
`include "AR_channel.sv"
`include "AW_channel.sv"
`include "R_channel.sv"
`include "W_channel.sv"
`include "B_channel.sv"
`include "Default_Slave.sv"
`include "Decoder.sv"
module AXI(
	input ACLK,
	input ARESETn,
    AXI_master_p.bridge master0,
    AXI_master_p.bridge master1,
    AXI_master_p.bridge master2,
    AXI_slave_p.bridge slave0,
    AXI_slave_p.bridge slave1,
    AXI_slave_p.bridge slave2,
    AXI_slave_p.bridge slave3,
    AXI_slave_p.bridge slave4,
    AXI_slave_p.bridge slave5
);
AXI_slave_p slave6();
logic [`AXI_MASTER_BITS-1:0] AW_Master;
logic [`AXI_SLAVE_BITS-1:0] AW_Slave;

Default_Slave default_slave(
    .clk(ACLK),
    .rst(ARESETn),
    .slave(slave6)
);

AR_channel AR_channel(
    .clk(ACLK),
    .rst(ARESETn),
	.ARID_M0   (master0.ARID),
	.ARADDR_M0 (master0.ARADDR),
	.ARLEN_M0  (master0.ARLEN),
	.ARSIZE_M0 (master0.ARSIZE),
	.ARBURST_M0(master0.ARBURST),
	.ARVALID_M0(master0.ARVALID),
    .ARREADY_M0(master0.ARREADY),
	.ARID_M1   (master1.ARID),
	.ARADDR_M1 (master1.ARADDR),
	.ARLEN_M1  (master1.ARLEN),
	.ARSIZE_M1 (master1.ARSIZE),
	.ARBURST_M1(master1.ARBURST),
	.ARVALID_M1(master1.ARVALID),
    .ARREADY_M1(master1.ARREADY),
	.ARID_M2   (master2.ARID),
	.ARADDR_M2 (master2.ARADDR),
	.ARLEN_M2  (master2.ARLEN),
	.ARSIZE_M2 (master2.ARSIZE),
	.ARBURST_M2(master2.ARBURST),
	.ARVALID_M2(master2.ARVALID),
    .ARREADY_M2(master2.ARREADY),
    .ARREADY_S0(slave0.ARREADY),
	.ARID_S0   (slave0.ARID   ),
	.ARADDR_S0 (slave0.ARADDR ),
	.ARLEN_S0  (slave0.ARLEN  ),
	.ARSIZE_S0 (slave0.ARSIZE ),
	.ARBURST_S0(slave0.ARBURST),
	.ARVALID_S0(slave0.ARVALID),
    .ARREADY_S1(slave1.ARREADY),
	.ARID_S1   (slave1.ARID   ),
	.ARADDR_S1 (slave1.ARADDR ),
	.ARLEN_S1  (slave1.ARLEN  ),
	.ARSIZE_S1 (slave1.ARSIZE ),
	.ARBURST_S1(slave1.ARBURST),
	.ARVALID_S1(slave1.ARVALID),
    .ARREADY_S2(slave2.ARREADY),
	.ARID_S2   (slave2.ARID   ),
	.ARADDR_S2 (slave2.ARADDR ),
	.ARLEN_S2  (slave2.ARLEN  ),
	.ARSIZE_S2 (slave2.ARSIZE ),
	.ARBURST_S2(slave2.ARBURST),
	.ARVALID_S2(slave2.ARVALID),
    .ARREADY_S3(slave3.ARREADY),
	.ARID_S3   (slave3.ARID   ),
	.ARADDR_S3 (slave3.ARADDR ),
	.ARLEN_S3  (slave3.ARLEN  ),
	.ARSIZE_S3 (slave3.ARSIZE ),
	.ARBURST_S3(slave3.ARBURST),
	.ARVALID_S3(slave3.ARVALID),
    .ARREADY_S4(slave4.ARREADY),
	.ARID_S4   (slave4.ARID   ),
	.ARADDR_S4 (slave4.ARADDR ),
	.ARLEN_S4  (slave4.ARLEN  ),
	.ARSIZE_S4 (slave4.ARSIZE ),
	.ARBURST_S4(slave4.ARBURST),
	.ARVALID_S4(slave4.ARVALID),
    .ARREADY_S5(slave5.ARREADY),
	.ARID_S5   (slave5.ARID   ),
	.ARADDR_S5 (slave5.ARADDR ),
	.ARLEN_S5  (slave5.ARLEN  ),
	.ARSIZE_S5 (slave5.ARSIZE ),
	.ARBURST_S5(slave5.ARBURST),
	.ARVALID_S5(slave5.ARVALID),
    .ARREADY_S6(slave6.ARREADY),
	.ARID_S6   (slave6.ARID   ),
	.ARADDR_S6 (slave6.ARADDR ),
	.ARLEN_S6  (slave6.ARLEN  ),
	.ARSIZE_S6 (slave6.ARSIZE ),
	.ARBURST_S6(slave6.ARBURST),
	.ARVALID_S6(slave6.ARVALID) 
);
AW_channel AW_channel(
    .clk(ACLK),
    .rst(ARESETn),
	.AWID_M0   (master0.AWID),
	.AWADDR_M0 (master0.AWADDR),
	.AWLEN_M0  (master0.AWLEN),
	.AWSIZE_M0 (master0.AWSIZE),
	.AWBURST_M0(master0.AWBURST),
	.AWVALID_M0(master0.AWVALID),
    .AWREADY_M0(master0.AWREADY),
	.AWID_M1   (master1.AWID),
	.AWADDR_M1 (master1.AWADDR),
	.AWLEN_M1  (master1.AWLEN),
	.AWSIZE_M1 (master1.AWSIZE),
	.AWBURST_M1(master1.AWBURST),
	.AWVALID_M1(master1.AWVALID),
    .AWREADY_M1(master1.AWREADY),
	.AWID_M2   (master2.AWID),
	.AWADDR_M2 (master2.AWADDR),
	.AWLEN_M2  (master2.AWLEN),
	.AWSIZE_M2 (master2.AWSIZE),
	.AWBURST_M2(master2.AWBURST),
	.AWVALID_M2(master2.AWVALID),
    .AWREADY_M2(master2.AWREADY),
    .AWREADY_S0(slave0.AWREADY),
	.AWID_S0   (slave0.AWID   ),
	.AWADDR_S0 (slave0.AWADDR ),
	.AWLEN_S0  (slave0.AWLEN  ),
	.AWSIZE_S0 (slave0.AWSIZE ),
	.AWBURST_S0(slave0.AWBURST),
	.AWVALID_S0(slave0.AWVALID),
    .AWREADY_S1(slave1.AWREADY),
	.AWID_S1   (slave1.AWID   ),
	.AWADDR_S1 (slave1.AWADDR ),
	.AWLEN_S1  (slave1.AWLEN  ),
	.AWSIZE_S1 (slave1.AWSIZE ),
	.AWBURST_S1(slave1.AWBURST),
	.AWVALID_S1(slave1.AWVALID),
    .AWREADY_S2(slave2.AWREADY),
	.AWID_S2   (slave2.AWID   ),
	.AWADDR_S2 (slave2.AWADDR ),
	.AWLEN_S2  (slave2.AWLEN  ),
	.AWSIZE_S2 (slave2.AWSIZE ),
	.AWBURST_S2(slave2.AWBURST),
	.AWVALID_S2(slave2.AWVALID),
    .AWREADY_S3(slave3.AWREADY),
	.AWID_S3   (slave3.AWID   ),
	.AWADDR_S3 (slave3.AWADDR ),
	.AWLEN_S3  (slave3.AWLEN  ),
	.AWSIZE_S3 (slave3.AWSIZE ),
	.AWBURST_S3(slave3.AWBURST),
	.AWVALID_S3(slave3.AWVALID),
    .AWREADY_S4(slave4.AWREADY),
	.AWID_S4   (slave4.AWID   ),
	.AWADDR_S4 (slave4.AWADDR ),
	.AWLEN_S4  (slave4.AWLEN  ),
	.AWSIZE_S4 (slave4.AWSIZE ),
	.AWBURST_S4(slave4.AWBURST),
	.AWVALID_S4(slave4.AWVALID),
    .AWREADY_S5(slave5.AWREADY),
	.AWID_S5   (slave5.AWID   ),
	.AWADDR_S5 (slave5.AWADDR ),
	.AWLEN_S5  (slave5.AWLEN  ),
	.AWSIZE_S5 (slave5.AWSIZE ),
	.AWBURST_S5(slave5.AWBURST),
	.AWVALID_S5(slave5.AWVALID),
    .AWREADY_S6(slave6.AWREADY),
	.AWID_S6   (slave6.AWID   ),
	.AWADDR_S6 (slave6.AWADDR ),
	.AWLEN_S6  (slave6.AWLEN  ),
	.AWSIZE_S6 (slave6.AWSIZE ),
	.AWBURST_S6(slave6.AWBURST),
	.AWVALID_S6(slave6.AWVALID),
    .Master(AW_Master),
    .slave(AW_Slave)
);

R_channel R_channel(
    .clk      (ACLK),
    .rst      (ARESETn),
    .RREADY_M0(master0.RREADY), 
	.RID_M0   (master0.RID   ),
	.RDATA_M0 (master0.RDATA ),
	.RRESP_M0 (master0.RRESP ),
	.RLAST_M0 (master0.RLAST ),
	.RVALID_M0(master0.RVALID),
    .RREADY_M1(master1.RREADY),
	.RID_M1   (master1.RID   ),
	.RDATA_M1 (master1.RDATA ),
	.RRESP_M1 (master1.RRESP ),
	.RLAST_M1 (master1.RLAST ),
	.RVALID_M1(master1.RVALID),
    .RREADY_M2(master2.RREADY),
	.RID_M2   (master2.RID   ),
	.RDATA_M2 (master2.RDATA ),
	.RRESP_M2 (master2.RRESP ),
	.RLAST_M2 (master2.RLAST ),
	.RVALID_M2(master2.RVALID),
	.RID_S0   (slave0.RID   ),
	.RDATA_S0 (slave0.RDATA ),
	.RRESP_S0 (slave0.RRESP ),
	.RLAST_S0 (slave0.RLAST ),
	.RVALID_S0(slave0.RVALID),
	.RREADY_S0(slave0.RREADY),
	.RID_S1   (slave1.RID   ),
	.RDATA_S1 (slave1.RDATA ),
	.RRESP_S1 (slave1.RRESP ),
	.RLAST_S1 (slave1.RLAST ),
	.RVALID_S1(slave1.RVALID),
	.RREADY_S1(slave1.RREADY),
	.RID_S2   (slave2.RID   ),
	.RDATA_S2 (slave2.RDATA ),
	.RRESP_S2 (slave2.RRESP ),
	.RLAST_S2 (slave2.RLAST ),
	.RVALID_S2(slave2.RVALID),
	.RREADY_S2(slave2.RREADY),
	.RID_S3   (slave3.RID   ),
	.RDATA_S3 (slave3.RDATA ),
	.RRESP_S3 (slave3.RRESP ),
	.RLAST_S3 (slave3.RLAST ),
	.RVALID_S3(slave3.RVALID),
	.RREADY_S3(slave3.RREADY),
	.RID_S4   (slave4.RID   ),
	.RDATA_S4 (slave4.RDATA ),
	.RRESP_S4 (slave4.RRESP ),
	.RLAST_S4 (slave4.RLAST ),
	.RVALID_S4(slave4.RVALID),
	.RREADY_S4(slave4.RREADY),
	.RID_S5   (slave5.RID   ),
	.RDATA_S5 (slave5.RDATA ),
	.RRESP_S5 (slave5.RRESP ),
	.RLAST_S5 (slave5.RLAST ),
	.RVALID_S5(slave5.RVALID),
	.RREADY_S5(slave5.RREADY),
	.RID_S6   (slave6.RID   ),
	.RDATA_S6 (slave6.RDATA ),
	.RRESP_S6 (slave6.RRESP ),
	.RLAST_S6 (slave6.RLAST ),
	.RVALID_S6(slave6.RVALID),
	.RREADY_S6(slave6.RREADY) 
);

W_channel w_channel(
    .clk       (ACLK),
    .rst       (ARESETn),
    .AW_slave  (AW_Slave),
	.WDATA_M0  (master0.WDATA  ),
	.WSTRB_M0  (master0.WSTRB  ),
	.WLAST_M0  (master0.WLAST  ),
	.WVALID_M0 (master0.WVALID ),
    .AWVALID_M0(master0.AWVALID),
	.WREADY_M0 (master0.WREADY ),
	.WDATA_M1  (master1.WDATA  ),
	.WSTRB_M1  (master1.WSTRB  ),
	.WLAST_M1  (master1.WLAST  ),
	.WVALID_M1 (master1.WVALID ),
    .AWVALID_M1(master1.AWVALID),
	.WREADY_M1 (master1.WREADY ),
	.WDATA_M2  (master2.WDATA  ),
	.WSTRB_M2  (master2.WSTRB  ),
	.WLAST_M2  (master2.WLAST  ),
	.WVALID_M2 (master2.WVALID ),
    .AWVALID_M2(master2.AWVALID),
	.WREADY_M2 (master2.WREADY ),
	.WDATA_S0  (slave0.WDATA   ),
	.WSTRB_S0  (slave0.WSTRB   ),
	.WLAST_S0  (slave0.WLAST   ),
	.WVALID_S0 (slave0.WVALID  ), 
	.WREADY_S0 (slave0.WREADY  ),
	.WDATA_S1  (slave1.WDATA   ),
	.WSTRB_S1  (slave1.WSTRB   ),
	.WLAST_S1  (slave1.WLAST   ),
	.WVALID_S1 (slave1.WVALID  ),
	.WREADY_S1 (slave1.WREADY  ),
	.WDATA_S2  (slave2.WDATA   ),
	.WSTRB_S2  (slave2.WSTRB   ),
	.WLAST_S2  (slave2.WLAST   ),
	.WVALID_S2 (slave2.WVALID  ),
	.WREADY_S2 (slave2.WREADY  ),
	.WDATA_S3  (slave3.WDATA   ),
	.WSTRB_S3  (slave3.WSTRB   ),
	.WLAST_S3  (slave3.WLAST   ),
	.WVALID_S3 (slave3.WVALID  ),
	.WREADY_S3 (slave3.WREADY  ),
	.WDATA_S4  (slave4.WDATA   ),
	.WSTRB_S4  (slave4.WSTRB   ),
	.WLAST_S4  (slave4.WLAST   ),
	.WVALID_S4 (slave4.WVALID  ),
	.WREADY_S4 (slave4.WREADY  ),
	.WDATA_S5  (slave5.WDATA   ),
	.WSTRB_S5  (slave5.WSTRB   ),
	.WLAST_S5  (slave5.WLAST   ),
	.WVALID_S5 (slave5.WVALID  ),
	.WREADY_S5 (slave5.WREADY  ),
	.WDATA_S6  (slave6.WDATA   ),
	.WSTRB_S6  (slave6.WSTRB   ),
	.WLAST_S6  (slave6.WLAST   ),
	.WVALID_S6 (slave6.WVALID  ),
	.WREADY_S6 (slave6.WREADY  ),
    .AWREADY_M0(master0.AWREADY),
    .AWREADY_M1(master1.AWREADY),
    .AWREADY_M2(master2.AWREADY)
);

B_channel B_channel(
    .clk(ACLK),
    .rst(ARESETn),
	.BID_M0   (master0.BID   ),
	.BRESP_M0 (master0.BRESP ),
	.BVALID_M0(master0.BVALID),
	.BREADY_M0(master0.BREADY),
	.BID_M1   (master1.BID   ),
	.BRESP_M1 (master1.BRESP ),
	.BVALID_M1(master1.BVALID),
	.BREADY_M1(master1.BREADY),
	.BID_M2   (master2.BID   ),
	.BRESP_M2 (master2.BRESP ),
	.BVALID_M2(master2.BVALID),
	.BREADY_M2(master2.BREADY),
	.BID_S0   (slave0.BID   ),
	.BRESP_S0 (slave0.BRESP ),
	.BVALID_S0(slave0.BVALID),
	.BREADY_S0(slave0.BREADY),
	.BID_S1   (slave1.BID   ),
	.BRESP_S1 (slave1.BRESP ),
	.BVALID_S1(slave1.BVALID),
	.BREADY_S1(slave1.BREADY),
    .BID_S2   (slave2.BID   ),
	.BRESP_S2 (slave2.BRESP ),
	.BVALID_S2(slave2.BVALID),
	.BREADY_S2(slave2.BREADY),
    .BID_S3   (slave3.BID   ),
	.BRESP_S3 (slave3.BRESP ),
	.BVALID_S3(slave3.BVALID),
	.BREADY_S3(slave3.BREADY),
    .BID_S4   (slave4.BID   ),
	.BRESP_S4 (slave4.BRESP ),
	.BVALID_S4(slave4.BVALID),
	.BREADY_S4(slave4.BREADY),
    .BID_S5   (slave5.BID   ),
	.BRESP_S5 (slave5.BRESP ),
	.BVALID_S5(slave5.BVALID),
	.BREADY_S5(slave5.BREADY),
	.BID_S6   (slave6.BID   ),
	.BRESP_S6 (slave6.BRESP ),
	.BVALID_S6(slave6.BVALID),
	.BREADY_S6(slave6.BREADY)
);
endmodule
