`include "AXI_define.svh"
module Arbiter(
    input clk,
    input rst,
    // Master0 interface
	input [`AXI_ID_BITS-1:0] ID_M0,
	input [`AXI_ADDR_BITS-1:0] ADDR_M0,
	input [`AXI_LEN_BITS-1:0] LEN_M0,
	input [`AXI_SIZE_BITS-1:0] SIZE_M0,
	input [1:0] BURST_M0,
	input VALID_M0,
    // Master1 interface
	input [`AXI_ID_BITS-1:0] ID_M1,
	input [`AXI_ADDR_BITS-1:0] ADDR_M1,
	input [`AXI_LEN_BITS-1:0] LEN_M1,
	input [`AXI_SIZE_BITS-1:0] SIZE_M1,
	input [1:0] BURST_M1,
	input VALID_M1,
    // Slave
    input READY,
    // output Master
	output logic [`AXI_IDS_BITS-1:0] ID_M,
	output logic [`AXI_ADDR_BITS-1:0] ADDR_M,
	output logic [`AXI_LEN_BITS-1:0] LEN_M,
	output logic [`AXI_SIZE_BITS-1:0] SIZE_M,
	output logic [1:0] BURST_M,
	output logic VALID_M,
    output logic READY_M0,
    output logic READY_M1,
	output logic [`AXI_MASTER_BITS-1:0] Master

);

logic LockM0;
logic LockM1;

always_ff@(posedge clk or negedge rst) begin
	if(~rst)begin
		LockM0 <= 1'b0;
		LockM1 <= 1'b0;
	end
	else begin
		LockM0 <= (LockM0 & READY) ? 1'b0 : (~VALID_M1 & VALID_M0 & ~READY) ? 1'b1 : LockM0;	
		LockM1 <= (LockM1 & READY) ? 1'b0 : (VALID_M1 & ~LockM0  & ~READY) ? 1'b1 : LockM1;	
	end
end

always_comb begin
	if((VALID_M1 & ~LockM0) | LockM1)
		Master = `AXI_MASTER1;
	else if (VALID_M0 | LockM0) 
		Master = `AXI_MASTER0;
	else 
		Master = `AXI_DEFAULT_MASTER;

end

always_comb begin
    case(Master)
        `AXI_MASTER0:begin
            ID_M = {`AXI_MASTER0,ID_M0};
            ADDR_M = ADDR_M0;
            LEN_M = LEN_M0;
            SIZE_M = SIZE_M0;
            BURST_M = BURST_M0;
            VALID_M = VALID_M0;
            READY_M0 = READY & VALID_M0;
            READY_M1 = 1'b0;
        end
        `AXI_MASTER1:begin
            ID_M = {`AXI_MASTER1,ID_M1};
            ADDR_M = ADDR_M1;
            LEN_M = LEN_M1;
            SIZE_M = SIZE_M1;
            BURST_M = BURST_M1;
            VALID_M = VALID_M1;
            READY_M0 = 1'b0;
            READY_M1 = READY & VALID_M1;
        end
        default:begin
            ID_M = {`AXI_DEFAULT_MASTER,`AXI_ID_BITS'b0};
            ADDR_M = `AXI_ADDR_BITS'b0;
            LEN_M = `AXI_LEN_BITS'b0;
            SIZE_M = `AXI_SIZE_BITS'b0;
            BURST_M = 2'b0;
            VALID_M = 1'b0;
            READY_M0 = 1'b0;
            READY_M1 = 1'b0;
        end
    endcase
end

endmodule
